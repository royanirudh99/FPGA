`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:57:42 06/24/2018 
// Design Name: 
// Module Name:    TX 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Transmiter( input CLK, input RST,input [7:0] DATA, output TX);
	reg [3:0] Count;	
	reg [10:0] IN = 11'b01001110001;			// 9600 Bauds at 12MHz			
	reg TX_register;
	wire Div_CLK;
	Clock_Divider CD1( CLK, IN,RST, Div_CLK);
	
	always @(posedge Div_CLK or posedge RST)
		begin
			if (RST)
				begin
					Count<=0;
					TX_register<=1;
				end
			else
				begin
					case (Count)
						4'b0000 : begin TX_register <= 0;Count<= Count +4'b0001; end
						4'b0001 : begin TX_register <= DATA[0];Count<= Count +4'b0001;end
						4'b0010 : begin TX_register <= DATA[1];Count<= Count +4'b0001;end
						4'b0011 : begin TX_register <= DATA[2];Count<= Count +4'b0001;end
						4'b0100 : begin TX_register <= DATA[3];Count<= Count +4'b0001;end
						4'b0101 : begin TX_register <= DATA[4];Count<= Count +4'b0001;end
						4'b0110 : begin TX_register <= DATA[5];Count<= Count +4'b0001;end
						4'b0111 : begin TX_register <= DATA[6];Count<= Count +4'b0001;end
						4'b1000 : begin TX_register <= DATA[7];Count<= Count +4'b0001;end
						4'b1001 : begin TX_register <= 1;Count<= Count +4'b0001;end					
						default : begin Count<=0; TX_register<=1; end
					endcase
				end
		end
		assign TX = TX_register;		
endmodule

